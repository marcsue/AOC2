library IEEE; 
use IEEE.STD_LOGIC_1164.all;

entity example410 is
port(
sw: in STD_LOGIC_VECTOR(4 downto 0);
ledG: out STD_LOGIC_VECTOR(3 downto 0));
end;
architecture synth of example410 is
begin
ledG <= sw(3 downto 0) when sw(4)= '1' else "ZZZZ";
end;